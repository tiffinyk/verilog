module bin2gry_test;
  parameter length = 4;
  //declare local variables
  reg [length-1:0] in ;
