module decode38(SW_In, LED_Out);
  input wire [2:0]SW_In;
  output wire [7:0]LED_Out;
endmodule
